/*******************************************************************************
    +-+-+-+-+-+-+-+-+-+-+ +-+-+-+-+-+-+-+-+-+-+-+-+ +-+-+ +-+-+-+-+-+-+-+-+
    |F|u|n|c|t|i|o|n|a|l| |V|e|r|i|f|i|c|a|t|i|o|n| |o|f| |H|a|r|d|w|a|r|e|
    +-+-+-+-+-+-+-+-+-+-+ +-+-+-+-+-+-+-+-+-+-+-+-+ +-+-+ +-+-+-+-+-+-+-+-+

    FILE            AXI_seq_lib.sv

    DESCRIPTION     includes all sequences

*******************************************************************************/


`include "sequences/AXILITE_base_seq.sv"
`include "sequences/AXIFULL_base_seq.sv"

`include "sequences/AXILITE_seq.sv"
`include "sequences/AXILITE2_seq.sv"
`include "sequences/AXIFULL_seq.sv"
`include "sequences/AXIFULL2_seq.sv"





